`include "global.v"

module speaker_control(

);


endmodule